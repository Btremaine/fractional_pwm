//////////////////////////////////////////////////////////////////////////////
// Module     : timescale.v                                                 //
// Description: This module contains the timescale for simulation.          //
//////////////////////////////////////////////////////////////////////////////

`timescale 1ns/1ps
