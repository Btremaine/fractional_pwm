//////////////////////////////////////////////////////////////////////////////
// Module     : defines.v                                                   //
// Description: This module contains system level definitions.              //
//////////////////////////////////////////////////////////////////////////////
`ifdef Veritak
`define BENCH
`else 
`undef BENCH
`endif
